`timescale 1ns/1ps
module Cgra6x6BlackBox(
            Config_Clock, 
            Config_Reset, 
            ConfigIn, 
            ConfigOut, 
            CGRA_Clock, 
            CGRA_Reset, 
            dataIn0,
            dataIn1,
            dataIn2,
            dataIn3,
            dataIn4,
            dataIn5,
            dataOut0,
            dataOut1,
            dataOut2,
            dataOut3,
            dataOut4,
            dataOut5,
            write,
            write_rq0,
            from_mem0,
            to_mem0,
            addr0,
            write_rq1,
            from_mem1,
            to_mem1,
            addr1,
            write_rq2,
            from_mem2,
            to_mem2,
            addr2,
            write_rq3,
            from_mem3,
            to_mem3,
            addr3,
            write_rq4,
            from_mem4,
            to_mem4,
            addr4,
            write_rq5,
            from_mem5,
            to_mem5,
            addr5);
    // Specifying the ports
    input Config_Clock, Config_Reset, ConfigIn;
    output ConfigOut;
    input CGRA_Clock, CGRA_Reset;

    output write_rq0;
    input [31:0] from_mem0;
    output [31:0] to_mem0;
    output [31:0] addr0;
    output write_rq1;
    input [31:0] from_mem1;
    output [31:0] to_mem1;
    output [31:0] addr1;
    output write_rq2;
    input [31:0] from_mem2;
    output [31:0] to_mem2;
    output [31:0] addr2;
    output write_rq3;
    input [31:0] from_mem3;
    output [31:0] to_mem3;
    output [31:0] addr3;
    output write_rq4;
    input [31:0] from_mem4;
    output [31:0] to_mem4;
    output [31:0] addr4;
    output write_rq5;
    input [31:0] from_mem5;
    output [31:0] to_mem5;
    output [31:0] addr5;

    wire [31:0] ext_io_top_0;
    wire [31:0] ext_io_top_1;
    wire [31:0] ext_io_top_2;
    wire [31:0] ext_io_top_3;
    wire [31:0] ext_io_top_4;
    wire [31:0] ext_io_top_5;

    input write;
    input [31:0] dataIn0;
    input [31:0] dataIn1;
    input [31:0] dataIn2;
    input [31:0] dataIn3;
    input [31:0] dataIn4;
    input [31:0] dataIn5;
    output [31:0] dataOut0;
    output [31:0] dataOut1;
    output [31:0] dataOut2;
    output [31:0] dataOut3;
    output [31:0] dataOut4;
    output [31:0] dataOut5;

    assign ext_io_top_0 = write? dataIn0 : 32'dz;
    assign ext_io_top_1 = write? dataIn1 : 32'dz;
    assign ext_io_top_2 = write? dataIn2 : 32'dz;
    assign ext_io_top_3 = write? dataIn3 : 32'dz;
    assign ext_io_top_4 = write? dataIn4 : 32'dz;
    assign ext_io_top_5 = write? dataIn5 : 32'dz;
    assign dataOut0 = ext_io_top_0;
    assign dataOut1 = ext_io_top_1;
    assign dataOut2 = ext_io_top_2;
    assign dataOut3 = ext_io_top_3;
    assign dataOut4 = ext_io_top_4;
    assign dataOut5 = ext_io_top_5;

    // Wires for the the config cells
    wire [2:0] DrfAddrIn0_sig;
    wire DrfAddrIn0_config;
    wire [2:0] DrfAddrIn1_sig;
    wire DrfAddrIn1_config;
    wire [2:0] DrfAddrIn2_sig;
    wire DrfAddrIn2_config;
    wire [2:0] DrfAddrIn3_sig;
    wire DrfAddrIn3_config;
    wire [2:0] DrfAddrIn4_sig;
    wire DrfAddrIn4_config;
    wire [2:0] DrfAddrIn5_sig;
    wire DrfAddrIn5_config;
    wire [2:0] DrfAddrOut0_sig;
    wire DrfAddrOut0_config;
    wire [2:0] DrfAddrOut1_sig;
    wire DrfAddrOut1_config;
    wire [2:0] DrfAddrOut10_sig;
    wire DrfAddrOut10_config;
    wire [2:0] DrfAddrOut11_sig;
    wire DrfAddrOut11_config;
    wire [2:0] DrfAddrOut2_sig;
    wire DrfAddrOut2_config;
    wire [2:0] DrfAddrOut3_sig;
    wire DrfAddrOut3_config;
    wire [2:0] DrfAddrOut4_sig;
    wire DrfAddrOut4_config;
    wire [2:0] DrfAddrOut5_sig;
    wire DrfAddrOut5_config;
    wire [2:0] DrfAddrOut6_sig;
    wire DrfAddrOut6_config;
    wire [2:0] DrfAddrOut7_sig;
    wire DrfAddrOut7_config;
    wire [2:0] DrfAddrOut8_sig;
    wire DrfAddrOut8_config;
    wire [2:0] DrfAddrOut9_sig;
    wire DrfAddrOut9_config;
    wire DrfWE0_sig;
    wire DrfWE0_config;
    wire DrfWE1_sig;
    wire DrfWE1_config;
    wire DrfWE2_sig;
    wire DrfWE2_config;
    wire DrfWE3_sig;
    wire DrfWE3_config;
    wire DrfWE4_sig;
    wire DrfWE4_config;
    wire DrfWE5_sig;
    wire DrfWE5_config;
    wire RfC0R1AddrIn0_sig;
    wire RfC0R1AddrIn0_config;
    wire RfC0R1AddrOut0_sig;
    wire RfC0R1AddrOut0_config;
    wire RfC0R1AddrOut1_sig;
    wire RfC0R1AddrOut1_config;
    wire RfC0R1WE_sig;
    wire RfC0R1WE_config;
    wire RfC0R2AddrIn0_sig;
    wire RfC0R2AddrIn0_config;
    wire RfC0R2AddrOut0_sig;
    wire RfC0R2AddrOut0_config;
    wire RfC0R2AddrOut1_sig;
    wire RfC0R2AddrOut1_config;
    wire RfC0R2WE_sig;
    wire RfC0R2WE_config;
    wire RfC0R3AddrIn0_sig;
    wire RfC0R3AddrIn0_config;
    wire RfC0R3AddrOut0_sig;
    wire RfC0R3AddrOut0_config;
    wire RfC0R3AddrOut1_sig;
    wire RfC0R3AddrOut1_config;
    wire RfC0R3WE_sig;
    wire RfC0R3WE_config;
    wire RfC0R4AddrIn0_sig;
    wire RfC0R4AddrIn0_config;
    wire RfC0R4AddrOut0_sig;
    wire RfC0R4AddrOut0_config;
    wire RfC0R4AddrOut1_sig;
    wire RfC0R4AddrOut1_config;
    wire RfC0R4WE_sig;
    wire RfC0R4WE_config;
    wire RfC0R5AddrIn0_sig;
    wire RfC0R5AddrIn0_config;
    wire RfC0R5AddrOut0_sig;
    wire RfC0R5AddrOut0_config;
    wire RfC0R5AddrOut1_sig;
    wire RfC0R5AddrOut1_config;
    wire RfC0R5WE_sig;
    wire RfC0R5WE_config;
    wire RfC1R1AddrIn0_sig;
    wire RfC1R1AddrIn0_config;
    wire RfC1R1AddrOut0_sig;
    wire RfC1R1AddrOut0_config;
    wire RfC1R1AddrOut1_sig;
    wire RfC1R1AddrOut1_config;
    wire RfC1R1WE_sig;
    wire RfC1R1WE_config;
    wire RfC1R2AddrIn0_sig;
    wire RfC1R2AddrIn0_config;
    wire RfC1R2AddrOut0_sig;
    wire RfC1R2AddrOut0_config;
    wire RfC1R2AddrOut1_sig;
    wire RfC1R2AddrOut1_config;
    wire RfC1R2WE_sig;
    wire RfC1R2WE_config;
    wire RfC1R3AddrIn0_sig;
    wire RfC1R3AddrIn0_config;
    wire RfC1R3AddrOut0_sig;
    wire RfC1R3AddrOut0_config;
    wire RfC1R3AddrOut1_sig;
    wire RfC1R3AddrOut1_config;
    wire RfC1R3WE_sig;
    wire RfC1R3WE_config;
    wire RfC1R4AddrIn0_sig;
    wire RfC1R4AddrIn0_config;
    wire RfC1R4AddrOut0_sig;
    wire RfC1R4AddrOut0_config;
    wire RfC1R4AddrOut1_sig;
    wire RfC1R4AddrOut1_config;
    wire RfC1R4WE_sig;
    wire RfC1R4WE_config;
    wire RfC1R5AddrIn0_sig;
    wire RfC1R5AddrIn0_config;
    wire RfC1R5AddrOut0_sig;
    wire RfC1R5AddrOut0_config;
    wire RfC1R5AddrOut1_sig;
    wire RfC1R5AddrOut1_config;
    wire RfC1R5WE_sig;
    wire RfC1R5WE_config;
    wire RfC2R1AddrIn0_sig;
    wire RfC2R1AddrIn0_config;
    wire RfC2R1AddrOut0_sig;
    wire RfC2R1AddrOut0_config;
    wire RfC2R1AddrOut1_sig;
    wire RfC2R1AddrOut1_config;
    wire RfC2R1WE_sig;
    wire RfC2R1WE_config;
    wire RfC2R2AddrIn0_sig;
    wire RfC2R2AddrIn0_config;
    wire RfC2R2AddrOut0_sig;
    wire RfC2R2AddrOut0_config;
    wire RfC2R2AddrOut1_sig;
    wire RfC2R2AddrOut1_config;
    wire RfC2R2WE_sig;
    wire RfC2R2WE_config;
    wire RfC2R3AddrIn0_sig;
    wire RfC2R3AddrIn0_config;
    wire RfC2R3AddrOut0_sig;
    wire RfC2R3AddrOut0_config;
    wire RfC2R3AddrOut1_sig;
    wire RfC2R3AddrOut1_config;
    wire RfC2R3WE_sig;
    wire RfC2R3WE_config;
    wire RfC2R4AddrIn0_sig;
    wire RfC2R4AddrIn0_config;
    wire RfC2R4AddrOut0_sig;
    wire RfC2R4AddrOut0_config;
    wire RfC2R4AddrOut1_sig;
    wire RfC2R4AddrOut1_config;
    wire RfC2R4WE_sig;
    wire RfC2R4WE_config;
    wire RfC2R5AddrIn0_sig;
    wire RfC2R5AddrIn0_config;
    wire RfC2R5AddrOut0_sig;
    wire RfC2R5AddrOut0_config;
    wire RfC2R5AddrOut1_sig;
    wire RfC2R5AddrOut1_config;
    wire RfC2R5WE_sig;
    wire RfC2R5WE_config;
    wire RfC3R1AddrIn0_sig;
    wire RfC3R1AddrIn0_config;
    wire RfC3R1AddrOut0_sig;
    wire RfC3R1AddrOut0_config;
    wire RfC3R1AddrOut1_sig;
    wire RfC3R1AddrOut1_config;
    wire RfC3R1WE_sig;
    wire RfC3R1WE_config;
    wire RfC3R2AddrIn0_sig;
    wire RfC3R2AddrIn0_config;
    wire RfC3R2AddrOut0_sig;
    wire RfC3R2AddrOut0_config;
    wire RfC3R2AddrOut1_sig;
    wire RfC3R2AddrOut1_config;
    wire RfC3R2WE_sig;
    wire RfC3R2WE_config;
    wire RfC3R3AddrIn0_sig;
    wire RfC3R3AddrIn0_config;
    wire RfC3R3AddrOut0_sig;
    wire RfC3R3AddrOut0_config;
    wire RfC3R3AddrOut1_sig;
    wire RfC3R3AddrOut1_config;
    wire RfC3R3WE_sig;
    wire RfC3R3WE_config;
    wire RfC3R4AddrIn0_sig;
    wire RfC3R4AddrIn0_config;
    wire RfC3R4AddrOut0_sig;
    wire RfC3R4AddrOut0_config;
    wire RfC3R4AddrOut1_sig;
    wire RfC3R4AddrOut1_config;
    wire RfC3R4WE_sig;
    wire RfC3R4WE_config;
    wire RfC3R5AddrIn0_sig;
    wire RfC3R5AddrIn0_config;
    wire RfC3R5AddrOut0_sig;
    wire RfC3R5AddrOut0_config;
    wire RfC3R5AddrOut1_sig;
    wire RfC3R5AddrOut1_config;
    wire RfC3R5WE_sig;
    wire RfC3R5WE_config;
    wire RfC4R1AddrIn0_sig;
    wire RfC4R1AddrIn0_config;
    wire RfC4R1AddrOut0_sig;
    wire RfC4R1AddrOut0_config;
    wire RfC4R1AddrOut1_sig;
    wire RfC4R1AddrOut1_config;
    wire RfC4R1WE_sig;
    wire RfC4R1WE_config;
    wire RfC4R2AddrIn0_sig;
    wire RfC4R2AddrIn0_config;
    wire RfC4R2AddrOut0_sig;
    wire RfC4R2AddrOut0_config;
    wire RfC4R2AddrOut1_sig;
    wire RfC4R2AddrOut1_config;
    wire RfC4R2WE_sig;
    wire RfC4R2WE_config;
    wire RfC4R3AddrIn0_sig;
    wire RfC4R3AddrIn0_config;
    wire RfC4R3AddrOut0_sig;
    wire RfC4R3AddrOut0_config;
    wire RfC4R3AddrOut1_sig;
    wire RfC4R3AddrOut1_config;
    wire RfC4R3WE_sig;
    wire RfC4R3WE_config;
    wire RfC4R4AddrIn0_sig;
    wire RfC4R4AddrIn0_config;
    wire RfC4R4AddrOut0_sig;
    wire RfC4R4AddrOut0_config;
    wire RfC4R4AddrOut1_sig;
    wire RfC4R4AddrOut1_config;
    wire RfC4R4WE_sig;
    wire RfC4R4WE_config;
    wire RfC4R5AddrIn0_sig;
    wire RfC4R5AddrIn0_config;
    wire RfC4R5AddrOut0_sig;
    wire RfC4R5AddrOut0_config;
    wire RfC4R5AddrOut1_sig;
    wire RfC4R5AddrOut1_config;
    wire RfC4R5WE_sig;
    wire RfC4R5WE_config;
    wire RfC5R1AddrIn0_sig;
    wire RfC5R1AddrIn0_config;
    wire RfC5R1AddrOut0_sig;
    wire RfC5R1AddrOut0_config;
    wire RfC5R1AddrOut1_sig;
    wire RfC5R1AddrOut1_config;
    wire RfC5R1WE_sig;
    wire RfC5R1WE_config;
    wire RfC5R2AddrIn0_sig;
    wire RfC5R2AddrIn0_config;
    wire RfC5R2AddrOut0_sig;
    wire RfC5R2AddrOut0_config;
    wire RfC5R2AddrOut1_sig;
    wire RfC5R2AddrOut1_config;
    wire RfC5R2WE_sig;
    wire RfC5R2WE_config;
    wire RfC5R3AddrIn0_sig;
    wire RfC5R3AddrIn0_config;
    wire RfC5R3AddrOut0_sig;
    wire RfC5R3AddrOut0_config;
    wire RfC5R3AddrOut1_sig;
    wire RfC5R3AddrOut1_config;
    wire RfC5R3WE_sig;
    wire RfC5R3WE_config;
    wire RfC5R4AddrIn0_sig;
    wire RfC5R4AddrIn0_config;
    wire RfC5R4AddrOut0_sig;
    wire RfC5R4AddrOut0_config;
    wire RfC5R4AddrOut1_sig;
    wire RfC5R4AddrOut1_config;
    wire RfC5R4WE_sig;
    wire RfC5R4WE_config;
    wire RfC5R5AddrIn0_sig;
    wire RfC5R5AddrIn0_config;
    wire RfC5R5AddrOut0_sig;
    wire RfC5R5AddrOut0_config;
    wire RfC5R5AddrOut1_sig;
    wire RfC5R5AddrOut1_config;
    wire RfC5R5WE_sig;
    wire RfC5R5WE_config;

    // Wires connecting the main module and submodules
    wire [31:0] io_top_1_out_sig;
    wire [31:0] io_top_2_out_sig;
    wire [31:0] io_top_0_out_sig;
    wire [31:0] io_top_3_out_sig;
    wire [31:0] io_top_4_out_sig;
    wire [31:0] io_top_5_out_sig;
    wire [31:0] mem_0_out_sig;
    wire [31:0] mem_1_out_sig;
    wire [31:0] mem_2_out_sig;
    wire [31:0] mem_3_out_sig;
    wire [31:0] mem_4_out_sig;
    wire [31:0] mem_5_out_sig;
    wire [31:0] pe_c0_r0_out_sig;
    wire [31:0] pe_c0_r0_fu_to_rf_sig;
    wire [31:0] pe_c0_r1_out_sig;
    wire [31:0] pe_c0_r1_fu_to_rf_sig;
    wire [31:0] pe_c0_r2_out_sig;
    wire [31:0] pe_c0_r2_fu_to_rf_sig;
    wire [31:0] pe_c0_r3_out_sig;
    wire [31:0] pe_c0_r3_fu_to_rf_sig;
    wire [31:0] pe_c0_r4_out_sig;
    wire [31:0] pe_c0_r4_fu_to_rf_sig;
    wire [31:0] pe_c0_r5_out_sig;
    wire [31:0] pe_c0_r5_fu_to_rf_sig;
    wire [31:0] pe_c1_r0_out_sig;
    wire [31:0] pe_c1_r0_fu_to_rf_sig;
    wire [31:0] pe_c1_r1_out_sig;
    wire [31:0] pe_c1_r1_fu_to_rf_sig;
    wire [31:0] pe_c1_r2_out_sig;
    wire [31:0] pe_c1_r2_fu_to_rf_sig;
    wire [31:0] pe_c1_r3_out_sig;
    wire [31:0] pe_c1_r3_fu_to_rf_sig;
    wire [31:0] pe_c1_r4_out_sig;
    wire [31:0] pe_c1_r4_fu_to_rf_sig;
    wire [31:0] pe_c1_r5_out_sig;
    wire [31:0] pe_c1_r5_fu_to_rf_sig;
    wire [31:0] pe_c2_r0_out_sig;
    wire [31:0] pe_c2_r0_fu_to_rf_sig;
    wire [31:0] pe_c2_r1_out_sig;
    wire [31:0] pe_c2_r1_fu_to_rf_sig;
    wire [31:0] pe_c2_r2_out_sig;
    wire [31:0] pe_c2_r2_fu_to_rf_sig;
    wire [31:0] pe_c2_r3_out_sig;
    wire [31:0] pe_c2_r3_fu_to_rf_sig;
    wire [31:0] pe_c2_r4_out_sig;
    wire [31:0] pe_c2_r4_fu_to_rf_sig;
    wire [31:0] pe_c2_r5_out_sig;
    wire [31:0] pe_c2_r5_fu_to_rf_sig;
    wire [31:0] pe_c3_r0_out_sig;
    wire [31:0] pe_c3_r0_fu_to_rf_sig;
    wire [31:0] pe_c3_r1_out_sig;
    wire [31:0] pe_c3_r1_fu_to_rf_sig;
    wire [31:0] pe_c3_r2_out_sig;
    wire [31:0] pe_c3_r2_fu_to_rf_sig;
    wire [31:0] pe_c3_r3_out_sig;
    wire [31:0] pe_c3_r3_fu_to_rf_sig;
    wire [31:0] pe_c3_r4_out_sig;
    wire [31:0] pe_c3_r4_fu_to_rf_sig;
    wire [31:0] pe_c3_r5_out_sig;
    wire [31:0] pe_c3_r5_fu_to_rf_sig;
    wire [31:0] pe_c4_r0_out_sig;
    wire [31:0] pe_c4_r0_fu_to_rf_sig;
    wire [31:0] pe_c4_r1_out_sig;
    wire [31:0] pe_c4_r1_fu_to_rf_sig;
    wire [31:0] pe_c4_r2_out_sig;
    wire [31:0] pe_c4_r2_fu_to_rf_sig;
    wire [31:0] pe_c4_r3_out_sig;
    wire [31:0] pe_c4_r3_fu_to_rf_sig;
    wire [31:0] pe_c4_r4_out_sig;
    wire [31:0] pe_c4_r4_fu_to_rf_sig;
    wire [31:0] pe_c4_r5_out_sig;
    wire [31:0] pe_c4_r5_fu_to_rf_sig;
    wire [31:0] pe_c5_r0_out_sig;
    wire [31:0] pe_c5_r0_fu_to_rf_sig;
    wire [31:0] pe_c5_r1_out_sig;
    wire [31:0] pe_c5_r1_fu_to_rf_sig;
    wire [31:0] pe_c5_r2_out_sig;
    wire [31:0] pe_c5_r2_fu_to_rf_sig;
    wire [31:0] pe_c5_r3_out_sig;
    wire [31:0] pe_c5_r3_fu_to_rf_sig;
    wire [31:0] pe_c5_r4_out_sig;
    wire [31:0] pe_c5_r4_fu_to_rf_sig;
    wire [31:0] pe_c5_r5_out_sig;
    wire [31:0] pe_c5_r5_fu_to_rf_sig;
    wire [31:0] drf_out0_sig;
    wire [31:0] drf_out1_sig;
    wire [31:0] drf_out2_sig;
    wire [31:0] drf_out3_sig;
    wire [31:0] drf_out4_sig;
    wire [31:0] drf_out5_sig;
    wire [31:0] drf_out6_sig;
    wire [31:0] drf_out7_sig;
    wire [31:0] drf_out8_sig;
    wire [31:0] drf_out9_sig;
    wire [31:0] drf_out10_sig;
    wire [31:0] drf_out11_sig;
    wire [31:0] rf_c0_r1_out0_sig;
    wire [31:0] rf_c0_r1_out1_sig;
    wire [31:0] rf_c0_r2_out0_sig;
    wire [31:0] rf_c0_r2_out1_sig;
    wire [31:0] rf_c0_r3_out0_sig;
    wire [31:0] rf_c0_r3_out1_sig;
    wire [31:0] rf_c0_r4_out0_sig;
    wire [31:0] rf_c0_r4_out1_sig;
    wire [31:0] rf_c0_r5_out0_sig;
    wire [31:0] rf_c0_r5_out1_sig;
    wire [31:0] rf_c1_r1_out0_sig;
    wire [31:0] rf_c1_r1_out1_sig;
    wire [31:0] rf_c1_r2_out0_sig;
    wire [31:0] rf_c1_r2_out1_sig;
    wire [31:0] rf_c1_r3_out0_sig;
    wire [31:0] rf_c1_r3_out1_sig;
    wire [31:0] rf_c1_r4_out0_sig;
    wire [31:0] rf_c1_r4_out1_sig;
    wire [31:0] rf_c1_r5_out0_sig;
    wire [31:0] rf_c1_r5_out1_sig;
    wire [31:0] rf_c2_r1_out0_sig;
    wire [31:0] rf_c2_r1_out1_sig;
    wire [31:0] rf_c2_r2_out0_sig;
    wire [31:0] rf_c2_r2_out1_sig;
    wire [31:0] rf_c2_r3_out0_sig;
    wire [31:0] rf_c2_r3_out1_sig;
    wire [31:0] rf_c2_r4_out0_sig;
    wire [31:0] rf_c2_r4_out1_sig;
    wire [31:0] rf_c2_r5_out0_sig;
    wire [31:0] rf_c2_r5_out1_sig;
    wire [31:0] rf_c3_r1_out0_sig;
    wire [31:0] rf_c3_r1_out1_sig;
    wire [31:0] rf_c3_r2_out0_sig;
    wire [31:0] rf_c3_r2_out1_sig;
    wire [31:0] rf_c3_r3_out0_sig;
    wire [31:0] rf_c3_r3_out1_sig;
    wire [31:0] rf_c3_r4_out0_sig;
    wire [31:0] rf_c3_r4_out1_sig;
    wire [31:0] rf_c3_r5_out0_sig;
    wire [31:0] rf_c3_r5_out1_sig;
    wire [31:0] rf_c4_r1_out0_sig;
    wire [31:0] rf_c4_r1_out1_sig;
    wire [31:0] rf_c4_r2_out0_sig;
    wire [31:0] rf_c4_r2_out1_sig;
    wire [31:0] rf_c4_r3_out0_sig;
    wire [31:0] rf_c4_r3_out1_sig;
    wire [31:0] rf_c4_r4_out0_sig;
    wire [31:0] rf_c4_r4_out1_sig;
    wire [31:0] rf_c4_r5_out0_sig;
    wire [31:0] rf_c4_r5_out1_sig;
    wire [31:0] rf_c5_r1_out0_sig;
    wire [31:0] rf_c5_r1_out1_sig;
    wire [31:0] rf_c5_r2_out0_sig;
    wire [31:0] rf_c5_r2_out1_sig;
    wire [31:0] rf_c5_r3_out0_sig;
    wire [31:0] rf_c5_r3_out1_sig;
    wire [31:0] rf_c5_r4_out0_sig;
    wire [31:0] rf_c5_r4_out1_sig;
    wire [31:0] rf_c5_r5_out0_sig;
    wire [31:0] rf_c5_r5_out1_sig;
    wire io_top_0_config;
    wire io_top_1_config;
    wire io_top_2_config;
    wire io_top_3_config;
    wire io_top_4_config;
    wire io_top_5_config;
    wire mem_0_config;
    wire mem_1_config;
    wire mem_2_config;
    wire mem_3_config;
    wire mem_4_config;
    wire mem_5_config;
    wire pe_c0_r0_config;
    wire pe_c0_r1_config;
    wire pe_c0_r2_config;
    wire pe_c0_r3_config;
    wire pe_c0_r4_config;
    wire pe_c0_r5_config;
    wire pe_c1_r0_config;
    wire pe_c1_r1_config;
    wire pe_c1_r2_config;
    wire pe_c1_r3_config;
    wire pe_c1_r4_config;
    wire pe_c1_r5_config;
    wire pe_c2_r0_config;
    wire pe_c2_r1_config;
    wire pe_c2_r2_config;
    wire pe_c2_r3_config;
    wire pe_c2_r4_config;
    wire pe_c2_r5_config;
    wire pe_c3_r0_config;
    wire pe_c3_r1_config;
    wire pe_c3_r2_config;
    wire pe_c3_r3_config;
    wire pe_c3_r4_config;
    wire pe_c3_r5_config;
    wire pe_c4_r0_config;
    wire pe_c4_r1_config;
    wire pe_c4_r2_config;
    wire pe_c4_r3_config;
    wire pe_c4_r4_config;
    wire pe_c4_r5_config;
    wire pe_c5_r0_config;
    wire pe_c5_r1_config;
    wire pe_c5_r2_config;
    wire pe_c5_r3_config;
    wire pe_c5_r4_config;
    wire pe_c5_r5_config;

    // Declaring the config cells
    ConfigCell #(3) DrfAddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(ConfigIn),
        .ConfigOut(DrfAddrIn0_config),
        .select(DrfAddrIn0_sig));
    ConfigCell #(3) DrfAddrIn1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn0_config),
        .ConfigOut(DrfAddrIn1_config),
        .select(DrfAddrIn1_sig));
    ConfigCell #(3) DrfAddrIn2 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn1_config),
        .ConfigOut(DrfAddrIn2_config),
        .select(DrfAddrIn2_sig));
    ConfigCell #(3) DrfAddrIn3 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn2_config),
        .ConfigOut(DrfAddrIn3_config),
        .select(DrfAddrIn3_sig));
    ConfigCell #(3) DrfAddrIn4 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn3_config),
        .ConfigOut(DrfAddrIn4_config),
        .select(DrfAddrIn4_sig));
    ConfigCell #(3) DrfAddrIn5 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn4_config),
        .ConfigOut(DrfAddrIn5_config),
        .select(DrfAddrIn5_sig));
    ConfigCell #(3) DrfAddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrIn5_config),
        .ConfigOut(DrfAddrOut0_config),
        .select(DrfAddrOut0_sig));
    ConfigCell #(3) DrfAddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut0_config),
        .ConfigOut(DrfAddrOut1_config),
        .select(DrfAddrOut1_sig));
    ConfigCell #(3) DrfAddrOut10 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut1_config),
        .ConfigOut(DrfAddrOut10_config),
        .select(DrfAddrOut10_sig));
    ConfigCell #(3) DrfAddrOut11 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut10_config),
        .ConfigOut(DrfAddrOut11_config),
        .select(DrfAddrOut11_sig));
    ConfigCell #(3) DrfAddrOut2 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut11_config),
        .ConfigOut(DrfAddrOut2_config),
        .select(DrfAddrOut2_sig));
    ConfigCell #(3) DrfAddrOut3 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut2_config),
        .ConfigOut(DrfAddrOut3_config),
        .select(DrfAddrOut3_sig));
    ConfigCell #(3) DrfAddrOut4 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut3_config),
        .ConfigOut(DrfAddrOut4_config),
        .select(DrfAddrOut4_sig));
    ConfigCell #(3) DrfAddrOut5 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut4_config),
        .ConfigOut(DrfAddrOut5_config),
        .select(DrfAddrOut5_sig));
    ConfigCell #(3) DrfAddrOut6 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut5_config),
        .ConfigOut(DrfAddrOut6_config),
        .select(DrfAddrOut6_sig));
    ConfigCell #(3) DrfAddrOut7 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut6_config),
        .ConfigOut(DrfAddrOut7_config),
        .select(DrfAddrOut7_sig));
    ConfigCell #(3) DrfAddrOut8 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut7_config),
        .ConfigOut(DrfAddrOut8_config),
        .select(DrfAddrOut8_sig));
    ConfigCell #(3) DrfAddrOut9 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut8_config),
        .ConfigOut(DrfAddrOut9_config),
        .select(DrfAddrOut9_sig));
    ConfigCell #(1) DrfWE0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfAddrOut9_config),
        .ConfigOut(DrfWE0_config),
        .select(DrfWE0_sig));
    ConfigCell #(1) DrfWE1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE0_config),
        .ConfigOut(DrfWE1_config),
        .select(DrfWE1_sig));
    ConfigCell #(1) DrfWE2 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE1_config),
        .ConfigOut(DrfWE2_config),
        .select(DrfWE2_sig));
    ConfigCell #(1) DrfWE3 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE2_config),
        .ConfigOut(DrfWE3_config),
        .select(DrfWE3_sig));
    ConfigCell #(1) DrfWE4 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE3_config),
        .ConfigOut(DrfWE4_config),
        .select(DrfWE4_sig));
    ConfigCell #(1) DrfWE5 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE4_config),
        .ConfigOut(DrfWE5_config),
        .select(DrfWE5_sig));
    ConfigCell #(1) RfC0R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(DrfWE5_config),
        .ConfigOut(RfC0R1AddrIn0_config),
        .select(RfC0R1AddrIn0_sig));
    ConfigCell #(1) RfC0R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R1AddrIn0_config),
        .ConfigOut(RfC0R1AddrOut0_config),
        .select(RfC0R1AddrOut0_sig));
    ConfigCell #(1) RfC0R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R1AddrOut0_config),
        .ConfigOut(RfC0R1AddrOut1_config),
        .select(RfC0R1AddrOut1_sig));
    ConfigCell #(1) RfC0R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R1AddrOut1_config),
        .ConfigOut(RfC0R1WE_config),
        .select(RfC0R1WE_sig));
    ConfigCell #(1) RfC0R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R1WE_config),
        .ConfigOut(RfC0R2AddrIn0_config),
        .select(RfC0R2AddrIn0_sig));
    ConfigCell #(1) RfC0R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R2AddrIn0_config),
        .ConfigOut(RfC0R2AddrOut0_config),
        .select(RfC0R2AddrOut0_sig));
    ConfigCell #(1) RfC0R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R2AddrOut0_config),
        .ConfigOut(RfC0R2AddrOut1_config),
        .select(RfC0R2AddrOut1_sig));
    ConfigCell #(1) RfC0R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R2AddrOut1_config),
        .ConfigOut(RfC0R2WE_config),
        .select(RfC0R2WE_sig));
    ConfigCell #(1) RfC0R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R2WE_config),
        .ConfigOut(RfC0R3AddrIn0_config),
        .select(RfC0R3AddrIn0_sig));
    ConfigCell #(1) RfC0R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R3AddrIn0_config),
        .ConfigOut(RfC0R3AddrOut0_config),
        .select(RfC0R3AddrOut0_sig));
    ConfigCell #(1) RfC0R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R3AddrOut0_config),
        .ConfigOut(RfC0R3AddrOut1_config),
        .select(RfC0R3AddrOut1_sig));
    ConfigCell #(1) RfC0R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R3AddrOut1_config),
        .ConfigOut(RfC0R3WE_config),
        .select(RfC0R3WE_sig));
    ConfigCell #(1) RfC0R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R3WE_config),
        .ConfigOut(RfC0R4AddrIn0_config),
        .select(RfC0R4AddrIn0_sig));
    ConfigCell #(1) RfC0R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R4AddrIn0_config),
        .ConfigOut(RfC0R4AddrOut0_config),
        .select(RfC0R4AddrOut0_sig));
    ConfigCell #(1) RfC0R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R4AddrOut0_config),
        .ConfigOut(RfC0R4AddrOut1_config),
        .select(RfC0R4AddrOut1_sig));
    ConfigCell #(1) RfC0R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R4AddrOut1_config),
        .ConfigOut(RfC0R4WE_config),
        .select(RfC0R4WE_sig));
    ConfigCell #(1) RfC0R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R4WE_config),
        .ConfigOut(RfC0R5AddrIn0_config),
        .select(RfC0R5AddrIn0_sig));
    ConfigCell #(1) RfC0R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R5AddrIn0_config),
        .ConfigOut(RfC0R5AddrOut0_config),
        .select(RfC0R5AddrOut0_sig));
    ConfigCell #(1) RfC0R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R5AddrOut0_config),
        .ConfigOut(RfC0R5AddrOut1_config),
        .select(RfC0R5AddrOut1_sig));
    ConfigCell #(1) RfC0R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R5AddrOut1_config),
        .ConfigOut(RfC0R5WE_config),
        .select(RfC0R5WE_sig));
    ConfigCell #(1) RfC1R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC0R5WE_config),
        .ConfigOut(RfC1R1AddrIn0_config),
        .select(RfC1R1AddrIn0_sig));
    ConfigCell #(1) RfC1R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R1AddrIn0_config),
        .ConfigOut(RfC1R1AddrOut0_config),
        .select(RfC1R1AddrOut0_sig));
    ConfigCell #(1) RfC1R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R1AddrOut0_config),
        .ConfigOut(RfC1R1AddrOut1_config),
        .select(RfC1R1AddrOut1_sig));
    ConfigCell #(1) RfC1R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R1AddrOut1_config),
        .ConfigOut(RfC1R1WE_config),
        .select(RfC1R1WE_sig));
    ConfigCell #(1) RfC1R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R1WE_config),
        .ConfigOut(RfC1R2AddrIn0_config),
        .select(RfC1R2AddrIn0_sig));
    ConfigCell #(1) RfC1R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R2AddrIn0_config),
        .ConfigOut(RfC1R2AddrOut0_config),
        .select(RfC1R2AddrOut0_sig));
    ConfigCell #(1) RfC1R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R2AddrOut0_config),
        .ConfigOut(RfC1R2AddrOut1_config),
        .select(RfC1R2AddrOut1_sig));
    ConfigCell #(1) RfC1R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R2AddrOut1_config),
        .ConfigOut(RfC1R2WE_config),
        .select(RfC1R2WE_sig));
    ConfigCell #(1) RfC1R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R2WE_config),
        .ConfigOut(RfC1R3AddrIn0_config),
        .select(RfC1R3AddrIn0_sig));
    ConfigCell #(1) RfC1R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R3AddrIn0_config),
        .ConfigOut(RfC1R3AddrOut0_config),
        .select(RfC1R3AddrOut0_sig));
    ConfigCell #(1) RfC1R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R3AddrOut0_config),
        .ConfigOut(RfC1R3AddrOut1_config),
        .select(RfC1R3AddrOut1_sig));
    ConfigCell #(1) RfC1R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R3AddrOut1_config),
        .ConfigOut(RfC1R3WE_config),
        .select(RfC1R3WE_sig));
    ConfigCell #(1) RfC1R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R3WE_config),
        .ConfigOut(RfC1R4AddrIn0_config),
        .select(RfC1R4AddrIn0_sig));
    ConfigCell #(1) RfC1R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R4AddrIn0_config),
        .ConfigOut(RfC1R4AddrOut0_config),
        .select(RfC1R4AddrOut0_sig));
    ConfigCell #(1) RfC1R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R4AddrOut0_config),
        .ConfigOut(RfC1R4AddrOut1_config),
        .select(RfC1R4AddrOut1_sig));
    ConfigCell #(1) RfC1R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R4AddrOut1_config),
        .ConfigOut(RfC1R4WE_config),
        .select(RfC1R4WE_sig));
    ConfigCell #(1) RfC1R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R4WE_config),
        .ConfigOut(RfC1R5AddrIn0_config),
        .select(RfC1R5AddrIn0_sig));
    ConfigCell #(1) RfC1R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R5AddrIn0_config),
        .ConfigOut(RfC1R5AddrOut0_config),
        .select(RfC1R5AddrOut0_sig));
    ConfigCell #(1) RfC1R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R5AddrOut0_config),
        .ConfigOut(RfC1R5AddrOut1_config),
        .select(RfC1R5AddrOut1_sig));
    ConfigCell #(1) RfC1R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R5AddrOut1_config),
        .ConfigOut(RfC1R5WE_config),
        .select(RfC1R5WE_sig));
    ConfigCell #(1) RfC2R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC1R5WE_config),
        .ConfigOut(RfC2R1AddrIn0_config),
        .select(RfC2R1AddrIn0_sig));
    ConfigCell #(1) RfC2R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R1AddrIn0_config),
        .ConfigOut(RfC2R1AddrOut0_config),
        .select(RfC2R1AddrOut0_sig));
    ConfigCell #(1) RfC2R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R1AddrOut0_config),
        .ConfigOut(RfC2R1AddrOut1_config),
        .select(RfC2R1AddrOut1_sig));
    ConfigCell #(1) RfC2R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R1AddrOut1_config),
        .ConfigOut(RfC2R1WE_config),
        .select(RfC2R1WE_sig));
    ConfigCell #(1) RfC2R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R1WE_config),
        .ConfigOut(RfC2R2AddrIn0_config),
        .select(RfC2R2AddrIn0_sig));
    ConfigCell #(1) RfC2R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R2AddrIn0_config),
        .ConfigOut(RfC2R2AddrOut0_config),
        .select(RfC2R2AddrOut0_sig));
    ConfigCell #(1) RfC2R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R2AddrOut0_config),
        .ConfigOut(RfC2R2AddrOut1_config),
        .select(RfC2R2AddrOut1_sig));
    ConfigCell #(1) RfC2R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R2AddrOut1_config),
        .ConfigOut(RfC2R2WE_config),
        .select(RfC2R2WE_sig));
    ConfigCell #(1) RfC2R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R2WE_config),
        .ConfigOut(RfC2R3AddrIn0_config),
        .select(RfC2R3AddrIn0_sig));
    ConfigCell #(1) RfC2R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R3AddrIn0_config),
        .ConfigOut(RfC2R3AddrOut0_config),
        .select(RfC2R3AddrOut0_sig));
    ConfigCell #(1) RfC2R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R3AddrOut0_config),
        .ConfigOut(RfC2R3AddrOut1_config),
        .select(RfC2R3AddrOut1_sig));
    ConfigCell #(1) RfC2R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R3AddrOut1_config),
        .ConfigOut(RfC2R3WE_config),
        .select(RfC2R3WE_sig));
    ConfigCell #(1) RfC2R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R3WE_config),
        .ConfigOut(RfC2R4AddrIn0_config),
        .select(RfC2R4AddrIn0_sig));
    ConfigCell #(1) RfC2R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R4AddrIn0_config),
        .ConfigOut(RfC2R4AddrOut0_config),
        .select(RfC2R4AddrOut0_sig));
    ConfigCell #(1) RfC2R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R4AddrOut0_config),
        .ConfigOut(RfC2R4AddrOut1_config),
        .select(RfC2R4AddrOut1_sig));
    ConfigCell #(1) RfC2R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R4AddrOut1_config),
        .ConfigOut(RfC2R4WE_config),
        .select(RfC2R4WE_sig));
    ConfigCell #(1) RfC2R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R4WE_config),
        .ConfigOut(RfC2R5AddrIn0_config),
        .select(RfC2R5AddrIn0_sig));
    ConfigCell #(1) RfC2R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R5AddrIn0_config),
        .ConfigOut(RfC2R5AddrOut0_config),
        .select(RfC2R5AddrOut0_sig));
    ConfigCell #(1) RfC2R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R5AddrOut0_config),
        .ConfigOut(RfC2R5AddrOut1_config),
        .select(RfC2R5AddrOut1_sig));
    ConfigCell #(1) RfC2R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R5AddrOut1_config),
        .ConfigOut(RfC2R5WE_config),
        .select(RfC2R5WE_sig));
    ConfigCell #(1) RfC3R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC2R5WE_config),
        .ConfigOut(RfC3R1AddrIn0_config),
        .select(RfC3R1AddrIn0_sig));
    ConfigCell #(1) RfC3R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R1AddrIn0_config),
        .ConfigOut(RfC3R1AddrOut0_config),
        .select(RfC3R1AddrOut0_sig));
    ConfigCell #(1) RfC3R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R1AddrOut0_config),
        .ConfigOut(RfC3R1AddrOut1_config),
        .select(RfC3R1AddrOut1_sig));
    ConfigCell #(1) RfC3R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R1AddrOut1_config),
        .ConfigOut(RfC3R1WE_config),
        .select(RfC3R1WE_sig));
    ConfigCell #(1) RfC3R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R1WE_config),
        .ConfigOut(RfC3R2AddrIn0_config),
        .select(RfC3R2AddrIn0_sig));
    ConfigCell #(1) RfC3R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R2AddrIn0_config),
        .ConfigOut(RfC3R2AddrOut0_config),
        .select(RfC3R2AddrOut0_sig));
    ConfigCell #(1) RfC3R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R2AddrOut0_config),
        .ConfigOut(RfC3R2AddrOut1_config),
        .select(RfC3R2AddrOut1_sig));
    ConfigCell #(1) RfC3R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R2AddrOut1_config),
        .ConfigOut(RfC3R2WE_config),
        .select(RfC3R2WE_sig));
    ConfigCell #(1) RfC3R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R2WE_config),
        .ConfigOut(RfC3R3AddrIn0_config),
        .select(RfC3R3AddrIn0_sig));
    ConfigCell #(1) RfC3R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R3AddrIn0_config),
        .ConfigOut(RfC3R3AddrOut0_config),
        .select(RfC3R3AddrOut0_sig));
    ConfigCell #(1) RfC3R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R3AddrOut0_config),
        .ConfigOut(RfC3R3AddrOut1_config),
        .select(RfC3R3AddrOut1_sig));
    ConfigCell #(1) RfC3R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R3AddrOut1_config),
        .ConfigOut(RfC3R3WE_config),
        .select(RfC3R3WE_sig));
    ConfigCell #(1) RfC3R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R3WE_config),
        .ConfigOut(RfC3R4AddrIn0_config),
        .select(RfC3R4AddrIn0_sig));
    ConfigCell #(1) RfC3R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R4AddrIn0_config),
        .ConfigOut(RfC3R4AddrOut0_config),
        .select(RfC3R4AddrOut0_sig));
    ConfigCell #(1) RfC3R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R4AddrOut0_config),
        .ConfigOut(RfC3R4AddrOut1_config),
        .select(RfC3R4AddrOut1_sig));
    ConfigCell #(1) RfC3R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R4AddrOut1_config),
        .ConfigOut(RfC3R4WE_config),
        .select(RfC3R4WE_sig));
    ConfigCell #(1) RfC3R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R4WE_config),
        .ConfigOut(RfC3R5AddrIn0_config),
        .select(RfC3R5AddrIn0_sig));
    ConfigCell #(1) RfC3R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R5AddrIn0_config),
        .ConfigOut(RfC3R5AddrOut0_config),
        .select(RfC3R5AddrOut0_sig));
    ConfigCell #(1) RfC3R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R5AddrOut0_config),
        .ConfigOut(RfC3R5AddrOut1_config),
        .select(RfC3R5AddrOut1_sig));
    ConfigCell #(1) RfC3R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R5AddrOut1_config),
        .ConfigOut(RfC3R5WE_config),
        .select(RfC3R5WE_sig));
    ConfigCell #(1) RfC4R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC3R5WE_config),
        .ConfigOut(RfC4R1AddrIn0_config),
        .select(RfC4R1AddrIn0_sig));
    ConfigCell #(1) RfC4R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R1AddrIn0_config),
        .ConfigOut(RfC4R1AddrOut0_config),
        .select(RfC4R1AddrOut0_sig));
    ConfigCell #(1) RfC4R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R1AddrOut0_config),
        .ConfigOut(RfC4R1AddrOut1_config),
        .select(RfC4R1AddrOut1_sig));
    ConfigCell #(1) RfC4R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R1AddrOut1_config),
        .ConfigOut(RfC4R1WE_config),
        .select(RfC4R1WE_sig));
    ConfigCell #(1) RfC4R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R1WE_config),
        .ConfigOut(RfC4R2AddrIn0_config),
        .select(RfC4R2AddrIn0_sig));
    ConfigCell #(1) RfC4R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R2AddrIn0_config),
        .ConfigOut(RfC4R2AddrOut0_config),
        .select(RfC4R2AddrOut0_sig));
    ConfigCell #(1) RfC4R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R2AddrOut0_config),
        .ConfigOut(RfC4R2AddrOut1_config),
        .select(RfC4R2AddrOut1_sig));
    ConfigCell #(1) RfC4R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R2AddrOut1_config),
        .ConfigOut(RfC4R2WE_config),
        .select(RfC4R2WE_sig));
    ConfigCell #(1) RfC4R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R2WE_config),
        .ConfigOut(RfC4R3AddrIn0_config),
        .select(RfC4R3AddrIn0_sig));
    ConfigCell #(1) RfC4R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R3AddrIn0_config),
        .ConfigOut(RfC4R3AddrOut0_config),
        .select(RfC4R3AddrOut0_sig));
    ConfigCell #(1) RfC4R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R3AddrOut0_config),
        .ConfigOut(RfC4R3AddrOut1_config),
        .select(RfC4R3AddrOut1_sig));
    ConfigCell #(1) RfC4R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R3AddrOut1_config),
        .ConfigOut(RfC4R3WE_config),
        .select(RfC4R3WE_sig));
    ConfigCell #(1) RfC4R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R3WE_config),
        .ConfigOut(RfC4R4AddrIn0_config),
        .select(RfC4R4AddrIn0_sig));
    ConfigCell #(1) RfC4R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R4AddrIn0_config),
        .ConfigOut(RfC4R4AddrOut0_config),
        .select(RfC4R4AddrOut0_sig));
    ConfigCell #(1) RfC4R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R4AddrOut0_config),
        .ConfigOut(RfC4R4AddrOut1_config),
        .select(RfC4R4AddrOut1_sig));
    ConfigCell #(1) RfC4R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R4AddrOut1_config),
        .ConfigOut(RfC4R4WE_config),
        .select(RfC4R4WE_sig));
    ConfigCell #(1) RfC4R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R4WE_config),
        .ConfigOut(RfC4R5AddrIn0_config),
        .select(RfC4R5AddrIn0_sig));
    ConfigCell #(1) RfC4R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R5AddrIn0_config),
        .ConfigOut(RfC4R5AddrOut0_config),
        .select(RfC4R5AddrOut0_sig));
    ConfigCell #(1) RfC4R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R5AddrOut0_config),
        .ConfigOut(RfC4R5AddrOut1_config),
        .select(RfC4R5AddrOut1_sig));
    ConfigCell #(1) RfC4R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R5AddrOut1_config),
        .ConfigOut(RfC4R5WE_config),
        .select(RfC4R5WE_sig));
    ConfigCell #(1) RfC5R1AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC4R5WE_config),
        .ConfigOut(RfC5R1AddrIn0_config),
        .select(RfC5R1AddrIn0_sig));
    ConfigCell #(1) RfC5R1AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R1AddrIn0_config),
        .ConfigOut(RfC5R1AddrOut0_config),
        .select(RfC5R1AddrOut0_sig));
    ConfigCell #(1) RfC5R1AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R1AddrOut0_config),
        .ConfigOut(RfC5R1AddrOut1_config),
        .select(RfC5R1AddrOut1_sig));
    ConfigCell #(1) RfC5R1WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R1AddrOut1_config),
        .ConfigOut(RfC5R1WE_config),
        .select(RfC5R1WE_sig));
    ConfigCell #(1) RfC5R2AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R1WE_config),
        .ConfigOut(RfC5R2AddrIn0_config),
        .select(RfC5R2AddrIn0_sig));
    ConfigCell #(1) RfC5R2AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R2AddrIn0_config),
        .ConfigOut(RfC5R2AddrOut0_config),
        .select(RfC5R2AddrOut0_sig));
    ConfigCell #(1) RfC5R2AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R2AddrOut0_config),
        .ConfigOut(RfC5R2AddrOut1_config),
        .select(RfC5R2AddrOut1_sig));
    ConfigCell #(1) RfC5R2WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R2AddrOut1_config),
        .ConfigOut(RfC5R2WE_config),
        .select(RfC5R2WE_sig));
    ConfigCell #(1) RfC5R3AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R2WE_config),
        .ConfigOut(RfC5R3AddrIn0_config),
        .select(RfC5R3AddrIn0_sig));
    ConfigCell #(1) RfC5R3AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R3AddrIn0_config),
        .ConfigOut(RfC5R3AddrOut0_config),
        .select(RfC5R3AddrOut0_sig));
    ConfigCell #(1) RfC5R3AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R3AddrOut0_config),
        .ConfigOut(RfC5R3AddrOut1_config),
        .select(RfC5R3AddrOut1_sig));
    ConfigCell #(1) RfC5R3WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R3AddrOut1_config),
        .ConfigOut(RfC5R3WE_config),
        .select(RfC5R3WE_sig));
    ConfigCell #(1) RfC5R4AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R3WE_config),
        .ConfigOut(RfC5R4AddrIn0_config),
        .select(RfC5R4AddrIn0_sig));
    ConfigCell #(1) RfC5R4AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R4AddrIn0_config),
        .ConfigOut(RfC5R4AddrOut0_config),
        .select(RfC5R4AddrOut0_sig));
    ConfigCell #(1) RfC5R4AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R4AddrOut0_config),
        .ConfigOut(RfC5R4AddrOut1_config),
        .select(RfC5R4AddrOut1_sig));
    ConfigCell #(1) RfC5R4WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R4AddrOut1_config),
        .ConfigOut(RfC5R4WE_config),
        .select(RfC5R4WE_sig));
    ConfigCell #(1) RfC5R5AddrIn0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R4WE_config),
        .ConfigOut(RfC5R5AddrIn0_config),
        .select(RfC5R5AddrIn0_sig));
    ConfigCell #(1) RfC5R5AddrOut0 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R5AddrIn0_config),
        .ConfigOut(RfC5R5AddrOut0_config),
        .select(RfC5R5AddrOut0_sig));
    ConfigCell #(1) RfC5R5AddrOut1 (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R5AddrOut0_config),
        .ConfigOut(RfC5R5AddrOut1_config),
        .select(RfC5R5AddrOut1_sig));
    ConfigCell #(1) RfC5R5WE (
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R5AddrOut1_config),
        .ConfigOut(RfC5R5WE_config),
        .select(RfC5R5WE_sig));

    // Declaring the submodules
    registerFile_6in_12out_32b #(3, 32) drf(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(DrfWE0_sig),
        .WE1(DrfWE1_sig),
        .WE2(DrfWE2_sig),
        .WE3(DrfWE3_sig),
        .WE4(DrfWE4_sig),
        .WE5(DrfWE5_sig),
        .address_in0(DrfAddrIn0_sig),
        .address_in1(DrfAddrIn1_sig),
        .address_in2(DrfAddrIn2_sig),
        .address_in3(DrfAddrIn3_sig),
        .address_in4(DrfAddrIn4_sig),
        .address_in5(DrfAddrIn5_sig),
        .address_out0(DrfAddrOut0_sig),
        .address_out1(DrfAddrOut1_sig),
        .address_out10(DrfAddrOut10_sig),
        .address_out11(DrfAddrOut11_sig),
        .address_out2(DrfAddrOut2_sig),
        .address_out3(DrfAddrOut3_sig),
        .address_out4(DrfAddrOut4_sig),
        .address_out5(DrfAddrOut5_sig),
        .address_out6(DrfAddrOut6_sig),
        .address_out7(DrfAddrOut7_sig),
        .address_out8(DrfAddrOut8_sig),
        .address_out9(DrfAddrOut9_sig),
        .in0(pe_c0_r0_fu_to_rf_sig),
        .in1(pe_c1_r0_fu_to_rf_sig),
        .in2(pe_c2_r0_fu_to_rf_sig),
        .in3(pe_c3_r0_fu_to_rf_sig),
        .in4(pe_c4_r0_fu_to_rf_sig),
        .in5(pe_c5_r0_fu_to_rf_sig),
        .out0(drf_out0_sig),
        .out1(drf_out1_sig),
        .out10(drf_out10_sig),
        .out11(drf_out11_sig),
        .out2(drf_out2_sig),
        .out3(drf_out3_sig),
        .out4(drf_out4_sig),
        .out5(drf_out5_sig),
        .out6(drf_out6_sig),
        .out7(drf_out7_sig),
        .out8(drf_out8_sig),
        .out9(drf_out9_sig));
    io_32b #(32) io_top_0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(RfC5R5WE_config),
        .ConfigOut(io_top_0_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_0),
        .in(pe_c0_r0_out_sig),
        .out(io_top_0_out_sig));
    io_32b #(32) io_top_1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_0_config),
        .ConfigOut(io_top_1_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_1),
        .in(pe_c1_r0_out_sig),
        .out(io_top_1_out_sig));
    io_32b #(32) io_top_2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_1_config),
        .ConfigOut(io_top_2_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_2),
        .in(pe_c2_r0_out_sig),
        .out(io_top_2_out_sig));
    io_32b #(32) io_top_3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_2_config),
        .ConfigOut(io_top_3_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_3),
        .in(pe_c3_r0_out_sig),
        .out(io_top_3_out_sig));
    io_32b #(32) io_top_4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_3_config),
        .ConfigOut(io_top_4_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_4),
        .in(pe_c4_r0_out_sig),
        .out(io_top_4_out_sig));
    io_32b #(32) io_top_5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_4_config),
        .ConfigOut(io_top_5_config),
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .bidir(ext_io_top_5),
        .in(pe_c5_r0_out_sig),
        .out(io_top_5_out_sig));
    memoryPort_6connect_32b mem_0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(io_top_5_config),
        .ConfigOut(mem_0_config),
        .in0(pe_c0_r0_out_sig),
        .in1(pe_c1_r0_out_sig),
        .in2(pe_c2_r0_out_sig),
        .in3(pe_c3_r0_out_sig),
        .in4(pe_c4_r0_out_sig),
        .in5(pe_c5_r0_out_sig),
        .out(mem_0_out_sig),
        .write_rq(write_rq0),
        .from_mem(from_mem0),
        .to_mem(to_mem0),
        .addr(addr0));
    memoryPort_6connect_32b mem_1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_0_config),
        .ConfigOut(mem_1_config),
        .in0(pe_c0_r1_out_sig),
        .in1(pe_c1_r1_out_sig),
        .in2(pe_c2_r1_out_sig),
        .in3(pe_c3_r1_out_sig),
        .in4(pe_c4_r1_out_sig),
        .in5(pe_c5_r1_out_sig),
        .out(mem_1_out_sig),
        .write_rq(write_rq1),
        .from_mem(from_mem1),
        .to_mem(to_mem1),
        .addr(addr1));
    memoryPort_6connect_32b mem_2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_1_config),
        .ConfigOut(mem_2_config),
        .in0(pe_c0_r2_out_sig),
        .in1(pe_c1_r2_out_sig),
        .in2(pe_c2_r2_out_sig),
        .in3(pe_c3_r2_out_sig),
        .in4(pe_c4_r2_out_sig),
        .in5(pe_c5_r2_out_sig),
        .out(mem_2_out_sig),
        .write_rq(write_rq2),
        .from_mem(from_mem2),
        .to_mem(to_mem2),
        .addr(addr2));
    memoryPort_6connect_32b mem_3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_2_config),
        .ConfigOut(mem_3_config),
        .in0(pe_c0_r3_out_sig),
        .in1(pe_c1_r3_out_sig),
        .in2(pe_c2_r3_out_sig),
        .in3(pe_c3_r3_out_sig),
        .in4(pe_c4_r3_out_sig),
        .in5(pe_c5_r3_out_sig),
        .out(mem_3_out_sig),
        .write_rq(write_rq3),
        .from_mem(from_mem3),
        .to_mem(to_mem3),
        .addr(addr3));
    memoryPort_6connect_32b mem_4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_3_config),
        .ConfigOut(mem_4_config),
        .in0(pe_c0_r4_out_sig),
        .in1(pe_c1_r4_out_sig),
        .in2(pe_c2_r4_out_sig),
        .in3(pe_c3_r4_out_sig),
        .in4(pe_c4_r4_out_sig),
        .in5(pe_c5_r4_out_sig),
        .out(mem_4_out_sig),
        .write_rq(write_rq4),
        .from_mem(from_mem4),
        .to_mem(to_mem4),
        .addr(addr4));
    memoryPort_6connect_32b mem_5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_4_config),
        .ConfigOut(mem_5_config),
        .in0(pe_c0_r5_out_sig),
        .in1(pe_c1_r5_out_sig),
        .in2(pe_c2_r5_out_sig),
        .in3(pe_c3_r5_out_sig),
        .in4(pe_c4_r5_out_sig),
        .in5(pe_c5_r5_out_sig),
        .out(mem_5_out_sig),
        .write_rq(write_rq5),
        .from_mem(from_mem5),
        .to_mem(to_mem5),
        .addr(addr5));
    adres_6in_vliw pe_c0_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(mem_5_config),
        .ConfigOut(pe_c0_r0_config),
        .fu_to_rf(pe_c0_r0_fu_to_rf_sig),
        .in0(io_top_0_out_sig),
        .in1(pe_c1_r0_out_sig),
        .in2(pe_c0_r1_out_sig),
        .in3(pe_c5_r0_out_sig),
        .in4(pe_c0_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c0_r0_out_sig),
        .rf_to_muxa(drf_out0_sig),
        .rf_to_muxout(drf_out1_sig));
    adres_5in_vliw pe_c0_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r0_config),
        .ConfigOut(pe_c0_r1_config),
        .fu_to_rf(pe_c0_r1_fu_to_rf_sig),
        .in0(pe_c0_r0_out_sig),
        .in1(pe_c1_r1_out_sig),
        .in2(pe_c0_r2_out_sig),
        .in3(pe_c5_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c0_r1_out_sig),
        .rf_to_muxa(rf_c0_r1_out0_sig),
        .rf_to_muxout(rf_c0_r1_out1_sig));
    adres_5in_vliw pe_c0_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r1_config),
        .ConfigOut(pe_c0_r2_config),
        .fu_to_rf(pe_c0_r2_fu_to_rf_sig),
        .in0(pe_c0_r1_out_sig),
        .in1(pe_c1_r2_out_sig),
        .in2(pe_c0_r3_out_sig),
        .in3(pe_c5_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c0_r2_out_sig),
        .rf_to_muxa(rf_c0_r2_out0_sig),
        .rf_to_muxout(rf_c0_r2_out1_sig));
    adres_5in_vliw pe_c0_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r2_config),
        .ConfigOut(pe_c0_r3_config),
        .fu_to_rf(pe_c0_r3_fu_to_rf_sig),
        .in0(pe_c0_r2_out_sig),
        .in1(pe_c1_r3_out_sig),
        .in2(pe_c0_r4_out_sig),
        .in3(pe_c5_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c0_r3_out_sig),
        .rf_to_muxa(rf_c0_r3_out0_sig),
        .rf_to_muxout(rf_c0_r3_out1_sig));
    adres_5in_vliw pe_c0_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r3_config),
        .ConfigOut(pe_c0_r4_config),
        .fu_to_rf(pe_c0_r4_fu_to_rf_sig),
        .in0(pe_c0_r3_out_sig),
        .in1(pe_c1_r4_out_sig),
        .in2(pe_c0_r5_out_sig),
        .in3(pe_c5_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c0_r4_out_sig),
        .rf_to_muxa(rf_c0_r4_out0_sig),
        .rf_to_muxout(rf_c0_r4_out1_sig));
    adres_5in_vliw pe_c0_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r4_config),
        .ConfigOut(pe_c0_r5_config),
        .fu_to_rf(pe_c0_r5_fu_to_rf_sig),
        .in0(pe_c0_r4_out_sig),
        .in1(pe_c1_r5_out_sig),
        .in2(pe_c0_r0_out_sig),
        .in3(pe_c5_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c0_r5_out_sig),
        .rf_to_muxa(rf_c0_r5_out0_sig),
        .rf_to_muxout(rf_c0_r5_out1_sig));
    adres_6in_vliw pe_c1_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c0_r5_config),
        .ConfigOut(pe_c1_r0_config),
        .fu_to_rf(pe_c1_r0_fu_to_rf_sig),
        .in0(io_top_1_out_sig),
        .in1(pe_c2_r0_out_sig),
        .in2(pe_c1_r1_out_sig),
        .in3(pe_c0_r0_out_sig),
        .in4(pe_c1_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c1_r0_out_sig),
        .rf_to_muxa(drf_out2_sig),
        .rf_to_muxout(drf_out3_sig));
    adres_5in_vliw pe_c1_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r0_config),
        .ConfigOut(pe_c1_r1_config),
        .fu_to_rf(pe_c1_r1_fu_to_rf_sig),
        .in0(pe_c1_r0_out_sig),
        .in1(pe_c2_r1_out_sig),
        .in2(pe_c1_r2_out_sig),
        .in3(pe_c0_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c1_r1_out_sig),
        .rf_to_muxa(rf_c1_r1_out0_sig),
        .rf_to_muxout(rf_c1_r1_out1_sig));
    adres_5in_vliw pe_c1_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r1_config),
        .ConfigOut(pe_c1_r2_config),
        .fu_to_rf(pe_c1_r2_fu_to_rf_sig),
        .in0(pe_c1_r1_out_sig),
        .in1(pe_c2_r2_out_sig),
        .in2(pe_c1_r3_out_sig),
        .in3(pe_c0_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c1_r2_out_sig),
        .rf_to_muxa(rf_c1_r2_out0_sig),
        .rf_to_muxout(rf_c1_r2_out1_sig));
    adres_5in_vliw pe_c1_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r2_config),
        .ConfigOut(pe_c1_r3_config),
        .fu_to_rf(pe_c1_r3_fu_to_rf_sig),
        .in0(pe_c1_r2_out_sig),
        .in1(pe_c2_r3_out_sig),
        .in2(pe_c1_r4_out_sig),
        .in3(pe_c0_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c1_r3_out_sig),
        .rf_to_muxa(rf_c1_r3_out0_sig),
        .rf_to_muxout(rf_c1_r3_out1_sig));
    adres_5in_vliw pe_c1_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r3_config),
        .ConfigOut(pe_c1_r4_config),
        .fu_to_rf(pe_c1_r4_fu_to_rf_sig),
        .in0(pe_c1_r3_out_sig),
        .in1(pe_c2_r4_out_sig),
        .in2(pe_c1_r5_out_sig),
        .in3(pe_c0_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c1_r4_out_sig),
        .rf_to_muxa(rf_c1_r4_out0_sig),
        .rf_to_muxout(rf_c1_r4_out1_sig));
    adres_5in_vliw pe_c1_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r4_config),
        .ConfigOut(pe_c1_r5_config),
        .fu_to_rf(pe_c1_r5_fu_to_rf_sig),
        .in0(pe_c1_r4_out_sig),
        .in1(pe_c2_r5_out_sig),
        .in2(pe_c1_r0_out_sig),
        .in3(pe_c0_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c1_r5_out_sig),
        .rf_to_muxa(rf_c1_r5_out0_sig),
        .rf_to_muxout(rf_c1_r5_out1_sig));
    adres_6in_vliw pe_c2_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c1_r5_config),
        .ConfigOut(pe_c2_r0_config),
        .fu_to_rf(pe_c2_r0_fu_to_rf_sig),
        .in0(io_top_2_out_sig),
        .in1(pe_c3_r0_out_sig),
        .in2(pe_c2_r1_out_sig),
        .in3(pe_c1_r0_out_sig),
        .in4(pe_c2_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c2_r0_out_sig),
        .rf_to_muxa(drf_out4_sig),
        .rf_to_muxout(drf_out5_sig));
    adres_5in_vliw pe_c2_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r0_config),
        .ConfigOut(pe_c2_r1_config),
        .fu_to_rf(pe_c2_r1_fu_to_rf_sig),
        .in0(pe_c2_r0_out_sig),
        .in1(pe_c3_r1_out_sig),
        .in2(pe_c2_r2_out_sig),
        .in3(pe_c1_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c2_r1_out_sig),
        .rf_to_muxa(rf_c2_r1_out0_sig),
        .rf_to_muxout(rf_c2_r1_out1_sig));
    adres_5in_vliw pe_c2_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r1_config),
        .ConfigOut(pe_c2_r2_config),
        .fu_to_rf(pe_c2_r2_fu_to_rf_sig),
        .in0(pe_c2_r1_out_sig),
        .in1(pe_c3_r2_out_sig),
        .in2(pe_c2_r3_out_sig),
        .in3(pe_c1_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c2_r2_out_sig),
        .rf_to_muxa(rf_c2_r2_out0_sig),
        .rf_to_muxout(rf_c2_r2_out1_sig));
    adres_5in_vliw pe_c2_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r2_config),
        .ConfigOut(pe_c2_r3_config),
        .fu_to_rf(pe_c2_r3_fu_to_rf_sig),
        .in0(pe_c2_r2_out_sig),
        .in1(pe_c3_r3_out_sig),
        .in2(pe_c2_r4_out_sig),
        .in3(pe_c1_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c2_r3_out_sig),
        .rf_to_muxa(rf_c2_r3_out0_sig),
        .rf_to_muxout(rf_c2_r3_out1_sig));
    adres_5in_vliw pe_c2_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r3_config),
        .ConfigOut(pe_c2_r4_config),
        .fu_to_rf(pe_c2_r4_fu_to_rf_sig),
        .in0(pe_c2_r3_out_sig),
        .in1(pe_c3_r4_out_sig),
        .in2(pe_c2_r5_out_sig),
        .in3(pe_c1_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c2_r4_out_sig),
        .rf_to_muxa(rf_c2_r4_out0_sig),
        .rf_to_muxout(rf_c2_r4_out1_sig));
    adres_5in_vliw pe_c2_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r4_config),
        .ConfigOut(pe_c2_r5_config),
        .fu_to_rf(pe_c2_r5_fu_to_rf_sig),
        .in0(pe_c2_r4_out_sig),
        .in1(pe_c3_r5_out_sig),
        .in2(pe_c2_r0_out_sig),
        .in3(pe_c1_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c2_r5_out_sig),
        .rf_to_muxa(rf_c2_r5_out0_sig),
        .rf_to_muxout(rf_c2_r5_out1_sig));
    adres_6in_vliw pe_c3_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c2_r5_config),
        .ConfigOut(pe_c3_r0_config),
        .fu_to_rf(pe_c3_r0_fu_to_rf_sig),
        .in0(io_top_3_out_sig),
        .in1(pe_c4_r0_out_sig),
        .in2(pe_c3_r1_out_sig),
        .in3(pe_c2_r0_out_sig),
        .in4(pe_c3_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c3_r0_out_sig),
        .rf_to_muxa(drf_out6_sig),
        .rf_to_muxout(drf_out7_sig));
    adres_5in_vliw pe_c3_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r0_config),
        .ConfigOut(pe_c3_r1_config),
        .fu_to_rf(pe_c3_r1_fu_to_rf_sig),
        .in0(pe_c3_r0_out_sig),
        .in1(pe_c4_r1_out_sig),
        .in2(pe_c3_r2_out_sig),
        .in3(pe_c2_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c3_r1_out_sig),
        .rf_to_muxa(rf_c3_r1_out0_sig),
        .rf_to_muxout(rf_c3_r1_out1_sig));
    adres_5in_vliw pe_c3_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r1_config),
        .ConfigOut(pe_c3_r2_config),
        .fu_to_rf(pe_c3_r2_fu_to_rf_sig),
        .in0(pe_c3_r1_out_sig),
        .in1(pe_c4_r2_out_sig),
        .in2(pe_c3_r3_out_sig),
        .in3(pe_c2_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c3_r2_out_sig),
        .rf_to_muxa(rf_c3_r2_out0_sig),
        .rf_to_muxout(rf_c3_r2_out1_sig));
    adres_5in_vliw pe_c3_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r2_config),
        .ConfigOut(pe_c3_r3_config),
        .fu_to_rf(pe_c3_r3_fu_to_rf_sig),
        .in0(pe_c3_r2_out_sig),
        .in1(pe_c4_r3_out_sig),
        .in2(pe_c3_r4_out_sig),
        .in3(pe_c2_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c3_r3_out_sig),
        .rf_to_muxa(rf_c3_r3_out0_sig),
        .rf_to_muxout(rf_c3_r3_out1_sig));
    adres_5in_vliw pe_c3_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r3_config),
        .ConfigOut(pe_c3_r4_config),
        .fu_to_rf(pe_c3_r4_fu_to_rf_sig),
        .in0(pe_c3_r3_out_sig),
        .in1(pe_c4_r4_out_sig),
        .in2(pe_c3_r5_out_sig),
        .in3(pe_c2_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c3_r4_out_sig),
        .rf_to_muxa(rf_c3_r4_out0_sig),
        .rf_to_muxout(rf_c3_r4_out1_sig));
    adres_5in_vliw pe_c3_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r4_config),
        .ConfigOut(pe_c3_r5_config),
        .fu_to_rf(pe_c3_r5_fu_to_rf_sig),
        .in0(pe_c3_r4_out_sig),
        .in1(pe_c4_r5_out_sig),
        .in2(pe_c3_r0_out_sig),
        .in3(pe_c2_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c3_r5_out_sig),
        .rf_to_muxa(rf_c3_r5_out0_sig),
        .rf_to_muxout(rf_c3_r5_out1_sig));
    adres_6in_vliw pe_c4_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c3_r5_config),
        .ConfigOut(pe_c4_r0_config),
        .fu_to_rf(pe_c4_r0_fu_to_rf_sig),
        .in0(io_top_4_out_sig),
        .in1(pe_c5_r0_out_sig),
        .in2(pe_c4_r1_out_sig),
        .in3(pe_c3_r0_out_sig),
        .in4(pe_c4_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c4_r0_out_sig),
        .rf_to_muxa(drf_out8_sig),
        .rf_to_muxout(drf_out9_sig));
    adres_5in_vliw pe_c4_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r0_config),
        .ConfigOut(pe_c4_r1_config),
        .fu_to_rf(pe_c4_r1_fu_to_rf_sig),
        .in0(pe_c4_r0_out_sig),
        .in1(pe_c5_r1_out_sig),
        .in2(pe_c4_r2_out_sig),
        .in3(pe_c3_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c4_r1_out_sig),
        .rf_to_muxa(rf_c4_r1_out0_sig),
        .rf_to_muxout(rf_c4_r1_out1_sig));
    adres_5in_vliw pe_c4_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r1_config),
        .ConfigOut(pe_c4_r2_config),
        .fu_to_rf(pe_c4_r2_fu_to_rf_sig),
        .in0(pe_c4_r1_out_sig),
        .in1(pe_c5_r2_out_sig),
        .in2(pe_c4_r3_out_sig),
        .in3(pe_c3_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c4_r2_out_sig),
        .rf_to_muxa(rf_c4_r2_out0_sig),
        .rf_to_muxout(rf_c4_r2_out1_sig));
    adres_5in_vliw pe_c4_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r2_config),
        .ConfigOut(pe_c4_r3_config),
        .fu_to_rf(pe_c4_r3_fu_to_rf_sig),
        .in0(pe_c4_r2_out_sig),
        .in1(pe_c5_r3_out_sig),
        .in2(pe_c4_r4_out_sig),
        .in3(pe_c3_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c4_r3_out_sig),
        .rf_to_muxa(rf_c4_r3_out0_sig),
        .rf_to_muxout(rf_c4_r3_out1_sig));
    adres_5in_vliw pe_c4_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r3_config),
        .ConfigOut(pe_c4_r4_config),
        .fu_to_rf(pe_c4_r4_fu_to_rf_sig),
        .in0(pe_c4_r3_out_sig),
        .in1(pe_c5_r4_out_sig),
        .in2(pe_c4_r5_out_sig),
        .in3(pe_c3_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c4_r4_out_sig),
        .rf_to_muxa(rf_c4_r4_out0_sig),
        .rf_to_muxout(rf_c4_r4_out1_sig));
    adres_5in_vliw pe_c4_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r4_config),
        .ConfigOut(pe_c4_r5_config),
        .fu_to_rf(pe_c4_r5_fu_to_rf_sig),
        .in0(pe_c4_r4_out_sig),
        .in1(pe_c5_r5_out_sig),
        .in2(pe_c4_r0_out_sig),
        .in3(pe_c3_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c4_r5_out_sig),
        .rf_to_muxa(rf_c4_r5_out0_sig),
        .rf_to_muxout(rf_c4_r5_out1_sig));
    adres_6in_vliw pe_c5_r0(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c4_r5_config),
        .ConfigOut(pe_c5_r0_config),
        .fu_to_rf(pe_c5_r0_fu_to_rf_sig),
        .in0(io_top_5_out_sig),
        .in1(pe_c0_r0_out_sig),
        .in2(pe_c5_r1_out_sig),
        .in3(pe_c4_r0_out_sig),
        .in4(pe_c5_r5_out_sig),
        .in5(mem_0_out_sig),
        .out(pe_c5_r0_out_sig),
        .rf_to_muxa(drf_out10_sig),
        .rf_to_muxout(drf_out11_sig));
    adres_5in_vliw pe_c5_r1(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c5_r0_config),
        .ConfigOut(pe_c5_r1_config),
        .fu_to_rf(pe_c5_r1_fu_to_rf_sig),
        .in0(pe_c5_r0_out_sig),
        .in1(pe_c0_r1_out_sig),
        .in2(pe_c5_r2_out_sig),
        .in3(pe_c4_r1_out_sig),
        .in4(mem_1_out_sig),
        .out(pe_c5_r1_out_sig),
        .rf_to_muxa(rf_c5_r1_out0_sig),
        .rf_to_muxout(rf_c5_r1_out1_sig));
    adres_5in_vliw pe_c5_r2(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c5_r1_config),
        .ConfigOut(pe_c5_r2_config),
        .fu_to_rf(pe_c5_r2_fu_to_rf_sig),
        .in0(pe_c5_r1_out_sig),
        .in1(pe_c0_r2_out_sig),
        .in2(pe_c5_r3_out_sig),
        .in3(pe_c4_r2_out_sig),
        .in4(mem_2_out_sig),
        .out(pe_c5_r2_out_sig),
        .rf_to_muxa(rf_c5_r2_out0_sig),
        .rf_to_muxout(rf_c5_r2_out1_sig));
    adres_5in_vliw pe_c5_r3(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c5_r2_config),
        .ConfigOut(pe_c5_r3_config),
        .fu_to_rf(pe_c5_r3_fu_to_rf_sig),
        .in0(pe_c5_r2_out_sig),
        .in1(pe_c0_r3_out_sig),
        .in2(pe_c5_r4_out_sig),
        .in3(pe_c4_r3_out_sig),
        .in4(mem_3_out_sig),
        .out(pe_c5_r3_out_sig),
        .rf_to_muxa(rf_c5_r3_out0_sig),
        .rf_to_muxout(rf_c5_r3_out1_sig));
    adres_5in_vliw pe_c5_r4(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c5_r3_config),
        .ConfigOut(pe_c5_r4_config),
        .fu_to_rf(pe_c5_r4_fu_to_rf_sig),
        .in0(pe_c5_r3_out_sig),
        .in1(pe_c0_r4_out_sig),
        .in2(pe_c5_r5_out_sig),
        .in3(pe_c4_r4_out_sig),
        .in4(mem_4_out_sig),
        .out(pe_c5_r4_out_sig),
        .rf_to_muxa(rf_c5_r4_out0_sig),
        .rf_to_muxout(rf_c5_r4_out1_sig));
    adres_5in_vliw pe_c5_r5(
        .Config_Clock(Config_Clock),
        .Config_Reset(Config_Reset),
        .ConfigIn(pe_c5_r4_config),
        .ConfigOut(pe_c5_r5_config),
        .fu_to_rf(pe_c5_r5_fu_to_rf_sig),
        .in0(pe_c5_r4_out_sig),
        .in1(pe_c0_r5_out_sig),
        .in2(pe_c5_r0_out_sig),
        .in3(pe_c4_r5_out_sig),
        .in4(mem_5_out_sig),
        .out(pe_c5_r5_out_sig),
        .rf_to_muxa(rf_c5_r5_out0_sig),
        .rf_to_muxout(rf_c5_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c0_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC0R1WE_sig),
        .address_in0(RfC0R1AddrIn0_sig),
        .address_out0(RfC0R1AddrOut0_sig),
        .address_out1(RfC0R1AddrOut1_sig),
        .in0(pe_c0_r1_fu_to_rf_sig),
        .out0(rf_c0_r1_out0_sig),
        .out1(rf_c0_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c0_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC0R2WE_sig),
        .address_in0(RfC0R2AddrIn0_sig),
        .address_out0(RfC0R2AddrOut0_sig),
        .address_out1(RfC0R2AddrOut1_sig),
        .in0(pe_c0_r2_fu_to_rf_sig),
        .out0(rf_c0_r2_out0_sig),
        .out1(rf_c0_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c0_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC0R3WE_sig),
        .address_in0(RfC0R3AddrIn0_sig),
        .address_out0(RfC0R3AddrOut0_sig),
        .address_out1(RfC0R3AddrOut1_sig),
        .in0(pe_c0_r3_fu_to_rf_sig),
        .out0(rf_c0_r3_out0_sig),
        .out1(rf_c0_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c0_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC0R4WE_sig),
        .address_in0(RfC0R4AddrIn0_sig),
        .address_out0(RfC0R4AddrOut0_sig),
        .address_out1(RfC0R4AddrOut1_sig),
        .in0(pe_c0_r4_fu_to_rf_sig),
        .out0(rf_c0_r4_out0_sig),
        .out1(rf_c0_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c0_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC0R5WE_sig),
        .address_in0(RfC0R5AddrIn0_sig),
        .address_out0(RfC0R5AddrOut0_sig),
        .address_out1(RfC0R5AddrOut1_sig),
        .in0(pe_c0_r5_fu_to_rf_sig),
        .out0(rf_c0_r5_out0_sig),
        .out1(rf_c0_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c1_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC1R1WE_sig),
        .address_in0(RfC1R1AddrIn0_sig),
        .address_out0(RfC1R1AddrOut0_sig),
        .address_out1(RfC1R1AddrOut1_sig),
        .in0(pe_c1_r1_fu_to_rf_sig),
        .out0(rf_c1_r1_out0_sig),
        .out1(rf_c1_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c1_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC1R2WE_sig),
        .address_in0(RfC1R2AddrIn0_sig),
        .address_out0(RfC1R2AddrOut0_sig),
        .address_out1(RfC1R2AddrOut1_sig),
        .in0(pe_c1_r2_fu_to_rf_sig),
        .out0(rf_c1_r2_out0_sig),
        .out1(rf_c1_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c1_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC1R3WE_sig),
        .address_in0(RfC1R3AddrIn0_sig),
        .address_out0(RfC1R3AddrOut0_sig),
        .address_out1(RfC1R3AddrOut1_sig),
        .in0(pe_c1_r3_fu_to_rf_sig),
        .out0(rf_c1_r3_out0_sig),
        .out1(rf_c1_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c1_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC1R4WE_sig),
        .address_in0(RfC1R4AddrIn0_sig),
        .address_out0(RfC1R4AddrOut0_sig),
        .address_out1(RfC1R4AddrOut1_sig),
        .in0(pe_c1_r4_fu_to_rf_sig),
        .out0(rf_c1_r4_out0_sig),
        .out1(rf_c1_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c1_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC1R5WE_sig),
        .address_in0(RfC1R5AddrIn0_sig),
        .address_out0(RfC1R5AddrOut0_sig),
        .address_out1(RfC1R5AddrOut1_sig),
        .in0(pe_c1_r5_fu_to_rf_sig),
        .out0(rf_c1_r5_out0_sig),
        .out1(rf_c1_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c2_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC2R1WE_sig),
        .address_in0(RfC2R1AddrIn0_sig),
        .address_out0(RfC2R1AddrOut0_sig),
        .address_out1(RfC2R1AddrOut1_sig),
        .in0(pe_c2_r1_fu_to_rf_sig),
        .out0(rf_c2_r1_out0_sig),
        .out1(rf_c2_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c2_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC2R2WE_sig),
        .address_in0(RfC2R2AddrIn0_sig),
        .address_out0(RfC2R2AddrOut0_sig),
        .address_out1(RfC2R2AddrOut1_sig),
        .in0(pe_c2_r2_fu_to_rf_sig),
        .out0(rf_c2_r2_out0_sig),
        .out1(rf_c2_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c2_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC2R3WE_sig),
        .address_in0(RfC2R3AddrIn0_sig),
        .address_out0(RfC2R3AddrOut0_sig),
        .address_out1(RfC2R3AddrOut1_sig),
        .in0(pe_c2_r3_fu_to_rf_sig),
        .out0(rf_c2_r3_out0_sig),
        .out1(rf_c2_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c2_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC2R4WE_sig),
        .address_in0(RfC2R4AddrIn0_sig),
        .address_out0(RfC2R4AddrOut0_sig),
        .address_out1(RfC2R4AddrOut1_sig),
        .in0(pe_c2_r4_fu_to_rf_sig),
        .out0(rf_c2_r4_out0_sig),
        .out1(rf_c2_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c2_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC2R5WE_sig),
        .address_in0(RfC2R5AddrIn0_sig),
        .address_out0(RfC2R5AddrOut0_sig),
        .address_out1(RfC2R5AddrOut1_sig),
        .in0(pe_c2_r5_fu_to_rf_sig),
        .out0(rf_c2_r5_out0_sig),
        .out1(rf_c2_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c3_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC3R1WE_sig),
        .address_in0(RfC3R1AddrIn0_sig),
        .address_out0(RfC3R1AddrOut0_sig),
        .address_out1(RfC3R1AddrOut1_sig),
        .in0(pe_c3_r1_fu_to_rf_sig),
        .out0(rf_c3_r1_out0_sig),
        .out1(rf_c3_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c3_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC3R2WE_sig),
        .address_in0(RfC3R2AddrIn0_sig),
        .address_out0(RfC3R2AddrOut0_sig),
        .address_out1(RfC3R2AddrOut1_sig),
        .in0(pe_c3_r2_fu_to_rf_sig),
        .out0(rf_c3_r2_out0_sig),
        .out1(rf_c3_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c3_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC3R3WE_sig),
        .address_in0(RfC3R3AddrIn0_sig),
        .address_out0(RfC3R3AddrOut0_sig),
        .address_out1(RfC3R3AddrOut1_sig),
        .in0(pe_c3_r3_fu_to_rf_sig),
        .out0(rf_c3_r3_out0_sig),
        .out1(rf_c3_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c3_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC3R4WE_sig),
        .address_in0(RfC3R4AddrIn0_sig),
        .address_out0(RfC3R4AddrOut0_sig),
        .address_out1(RfC3R4AddrOut1_sig),
        .in0(pe_c3_r4_fu_to_rf_sig),
        .out0(rf_c3_r4_out0_sig),
        .out1(rf_c3_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c3_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC3R5WE_sig),
        .address_in0(RfC3R5AddrIn0_sig),
        .address_out0(RfC3R5AddrOut0_sig),
        .address_out1(RfC3R5AddrOut1_sig),
        .in0(pe_c3_r5_fu_to_rf_sig),
        .out0(rf_c3_r5_out0_sig),
        .out1(rf_c3_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c4_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC4R1WE_sig),
        .address_in0(RfC4R1AddrIn0_sig),
        .address_out0(RfC4R1AddrOut0_sig),
        .address_out1(RfC4R1AddrOut1_sig),
        .in0(pe_c4_r1_fu_to_rf_sig),
        .out0(rf_c4_r1_out0_sig),
        .out1(rf_c4_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c4_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC4R2WE_sig),
        .address_in0(RfC4R2AddrIn0_sig),
        .address_out0(RfC4R2AddrOut0_sig),
        .address_out1(RfC4R2AddrOut1_sig),
        .in0(pe_c4_r2_fu_to_rf_sig),
        .out0(rf_c4_r2_out0_sig),
        .out1(rf_c4_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c4_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC4R3WE_sig),
        .address_in0(RfC4R3AddrIn0_sig),
        .address_out0(RfC4R3AddrOut0_sig),
        .address_out1(RfC4R3AddrOut1_sig),
        .in0(pe_c4_r3_fu_to_rf_sig),
        .out0(rf_c4_r3_out0_sig),
        .out1(rf_c4_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c4_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC4R4WE_sig),
        .address_in0(RfC4R4AddrIn0_sig),
        .address_out0(RfC4R4AddrOut0_sig),
        .address_out1(RfC4R4AddrOut1_sig),
        .in0(pe_c4_r4_fu_to_rf_sig),
        .out0(rf_c4_r4_out0_sig),
        .out1(rf_c4_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c4_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC4R5WE_sig),
        .address_in0(RfC4R5AddrIn0_sig),
        .address_out0(RfC4R5AddrOut0_sig),
        .address_out1(RfC4R5AddrOut1_sig),
        .in0(pe_c4_r5_fu_to_rf_sig),
        .out0(rf_c4_r5_out0_sig),
        .out1(rf_c4_r5_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c5_r1(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC5R1WE_sig),
        .address_in0(RfC5R1AddrIn0_sig),
        .address_out0(RfC5R1AddrOut0_sig),
        .address_out1(RfC5R1AddrOut1_sig),
        .in0(pe_c5_r1_fu_to_rf_sig),
        .out0(rf_c5_r1_out0_sig),
        .out1(rf_c5_r1_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c5_r2(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC5R2WE_sig),
        .address_in0(RfC5R2AddrIn0_sig),
        .address_out0(RfC5R2AddrOut0_sig),
        .address_out1(RfC5R2AddrOut1_sig),
        .in0(pe_c5_r2_fu_to_rf_sig),
        .out0(rf_c5_r2_out0_sig),
        .out1(rf_c5_r2_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c5_r3(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC5R3WE_sig),
        .address_in0(RfC5R3AddrIn0_sig),
        .address_out0(RfC5R3AddrOut0_sig),
        .address_out1(RfC5R3AddrOut1_sig),
        .in0(pe_c5_r3_fu_to_rf_sig),
        .out0(rf_c5_r3_out0_sig),
        .out1(rf_c5_r3_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c5_r4(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC5R4WE_sig),
        .address_in0(RfC5R4AddrIn0_sig),
        .address_out0(RfC5R4AddrOut0_sig),
        .address_out1(RfC5R4AddrOut1_sig),
        .in0(pe_c5_r4_fu_to_rf_sig),
        .out0(rf_c5_r4_out0_sig),
        .out1(rf_c5_r4_out1_sig));
    registerFile_1in_2out_32b #(1, 32) rf_c5_r5(
        .CGRA_Clock(CGRA_Clock),
        .CGRA_Reset(CGRA_Reset),
        .WE0(RfC5R5WE_sig),
        .address_in0(RfC5R5AddrIn0_sig),
        .address_out0(RfC5R5AddrOut0_sig),
        .address_out1(RfC5R5AddrOut1_sig),
        .in0(pe_c5_r5_fu_to_rf_sig),
        .out0(rf_c5_r5_out0_sig),
        .out1(rf_c5_r5_out1_sig));
    assign ConfigOut = pe_c5_r5_config;
endmodule

